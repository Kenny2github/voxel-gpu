module pixel_shader #(
    parameter ROW = 0,
    parameter COL = 0,
    parameter ROW_BITS = 8,
    parameter COL_BITS = 8,
    parameter COORD_BITS = 8,
    parameter PALETTE_BITS = 8,
    parameter FRAC_BITS = 8,
    parameter PIXEL_BITS = 8
) (
    input logic do_rasterize,
    input logic do_shade,
    input logic [COORD_BITS-1:0] voxel_x,
    input logic [COORD_BITS-1:0] voxel_y,
    input logic [COORD_BITS-1:0] voxel_z,
    input logic [PALETTE_BITS-1:0] voxel_id,
    input logic signed [COORD_BITS+FRAC_BITS-1:0] cam_pos_x,
    input logic signed [COORD_BITS+FRAC_BITS-1:0] cam_pos_y,
    input logic signed [COORD_BITS+FRAC_BITS-1:0] cam_pos_z,
    input logic signed [COORD_BITS+FRAC_BITS-1:0] cam_look_x,
    input logic signed [COORD_BITS+FRAC_BITS-1:0] cam_look_y,
    input logic signed [COORD_BITS+FRAC_BITS-1:0] cam_look_z,
    input logic [ROW_BITS-1:0] row,
    input logic [COL_BITS-1:0] col,
    output logic rasterizing_done,
    output logic shading_done,
    output wire [PIXEL_BITS-1:0] pixel,
    input logic reset,
    input logic clock
);
  enum logic [3:0] {
    IDLE,
    MEASURE,
    STORE_VOXEL,
    DONE_RASTERIZING,
    STORE_PIXEL,
    DONE_SHADING
  }
      state, next_state;

  logic [PIXEL_BITS-1:0] _pixel;
  assign pixel = (row == ROW && col == COL) ? _pixel : 'z;

  logic [COORD_BITS+FRAC_BITS-1:0] tAx, tAy, tAz, tBx, tBy, tBz;

  assign tAx = {({voxel_x, FRAC_BITS'(0)} - cam_pos_x), FRAC_BITS'(0)} / (cam_look_x || 1);
  assign tAy = {({voxel_y, FRAC_BITS'(0)} - cam_pos_y), FRAC_BITS'(0)} / (cam_look_y || 1);
  assign tAz = {({voxel_z, FRAC_BITS'(0)} - cam_pos_z), FRAC_BITS'(0)} / (cam_look_z || 1);
  assign tBx = {({voxel_x + 1'b1, FRAC_BITS'(0)} - cam_pos_x), FRAC_BITS'(0)} / (cam_look_x || 1);
  assign tBy = {({voxel_y + 1'b1, FRAC_BITS'(0)} - cam_pos_y), FRAC_BITS'(0)} / (cam_look_y || 1);
  assign tBz = {({voxel_z + 1'b1, FRAC_BITS'(0)} - cam_pos_z), FRAC_BITS'(0)} / (cam_look_z || 1);

  always_ff @(posedge clock, posedge reset) begin
    if (reset) begin
      state <= IDLE;
    end else begin
      state <= next_state;
    end
  end

  always_comb begin
    case (state)
      IDLE: begin
        if (do_rasterize) next_state = MEASURE;
        else if (do_shade) next_state = STORE_PIXEL;
        else next_state = IDLE;
      end
      MEASURE: begin
        next_state = STORE_VOXEL;
      end
      STORE_VOXEL: begin
        next_state = DONE_RASTERIZING;
      end
      DONE_RASTERIZING: begin
        if (do_rasterize) next_state = MEASURE;
        else next_state = IDLE;
      end
      STORE_PIXEL: begin
        next_state = DONE_SHADING;
      end
      DONE_SHADING: begin
        if (do_shade) next_state = STORE_PIXEL;
        else next_state = IDLE;
      end
    endcase
  end

endmodule
